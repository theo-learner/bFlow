module test(A, B, out); 
	input A;
	input B;
	output out;

	assign out = A & B;  
endmodule
