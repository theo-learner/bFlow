/*	File:	decode.v	  						*/

/*	module name: decode						*/

/*	Description: decode */

/*		Perform 24 bit logical operations	*/


/*==============================================================================*/


/********************************************************************************/
/*																				*/
/*	module:																		*/
/*																				*/
/********************************************************************************/

module decode (
	in,
	out
	);


/*============	I/O direction	================================================*/

input [4:0] 	in;
output [`databus]	out;

/*==============================================================================*/



/*============		I/O type	================================================*/

wire [`databus]	 out;

/*==============================================================================*/


/*===========	Function Declarations	========================================*/


/*--------------------------------------------------------------------------------------*/
/*																						*/
/*	function:	power_of_2																*/
/*																						*/
/*	Calculates 2 ^ -(power), where n is a 5 bit number											*/
/*																						*/
/*--------------------------------------------------------------------------------------*/

function [24:0] power_of_2;

input [4:0] power;	/* The register to be tested */ 

begin
	case (power)
			5'b00001	:	power_of_2 = 24'h400000;
			5'b00010	:	power_of_2 = 24'h200000;
			5'b00011	:	power_of_2 = 24'h100000;
			5'b00100	:	power_of_2 = 24'h080000;
			5'b00101	:	power_of_2 = 24'h040000;
			5'b00110	:	power_of_2 = 24'h020000;
			5'b00111	:	power_of_2 = 24'h010000;
			5'b01000	:	power_of_2 = 24'h008000;
			5'b01001	:	power_of_2 = 24'h004000;
			5'b01010	:	power_of_2 = 24'h002000;
			5'b01011	:	power_of_2 = 24'h001000;
			5'b01100	:	power_of_2 = 24'h000800;
			5'b01101	:	power_of_2 = 24'h000400;
			5'b01110	:	power_of_2 = 24'h000200;
			5'b01111	:	power_of_2 = 24'h000100;
			5'b10000	:	power_of_2 = 24'h000080;
			5'b10001	:	power_of_2 = 24'h000040;
			5'b10010	:	power_of_2 = 24'h000020;
			5'b10011	:	power_of_2 = 24'h000010;
			5'b10100	:	power_of_2 = 24'h000008;
			5'b10101	:	power_of_2 = 24'h000004;
			5'b10110	:	power_of_2 = 24'h000002;
			5'b10111	:	power_of_2 = 24'h000001;
			default		:	/* ILLEGAL, set to 0 */
							power_of_2 = 24'h000000;
	endcase		/* power */
end
endfunction /* power_of_2 */



/*==============================================================================*/
/*	processes																	*/
/*==============================================================================*/

assign out =  power_of_2(in);


endmodule	/* end module */
