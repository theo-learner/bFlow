/*	File:	core.v	  						*/

/*	module name: core						*/

/*	Description: The Motorola 56K core module - comprises of the following units:	*/
/*				 agu 			The address generation unit							*/
/*				 data_alu		The data ALU										*/
/*				 bus_switch		The internal data bus switch						*/
/*				 pcu			The program control unit							*/

/*	Author: Nitzan Weineberg */

/*==============================================================================*/


/********************************************************************************/
/*																				*/
/*	module:	core1																*/
/*																				*/
/********************************************************************************/

module cmudsp(
	reset,
	PDB,
	XDB,
	YDB,
	PAB,
	XAB,
	XWRITE,
	XREAD,
	YAB,
	YWRITE,
	YREAD,
	Clk
	);


/*============	I/O direction	================================================*/

input reset;
input [`databus] PDB;
inout [`databus] XDB;
inout [`databus] YDB;

output [`addrbus] PAB;

output [`addrbus] XAB;
output XWRITE;
output XREAD;

output [`addrbus] YAB;
output YWRITE;
output YREAD;

input Clk;

/*==============================================================================*/



/*============		I/O type	================================================*/
wire reset;
wire [`databus] PDB;
wire [`databus] XDB;
wire [`databus] YDB;

wor [`addrbus] PAB;

wire [`addrbus] XAB;
wire XWRITE;
wire XREAD;

wire [`addrbus] YAB;
wire YWRITE;
wire YREAD;

wire Clk;

/*==============================================================================*/



/*===========	Internal Nets	================================================*/

wire [`databus] GDB;		/* the GDB 24-bit internal bi-directional data bus */

wire [`addrbus] GDB_PCU;	/* GDB connection to the PCU but is 16-bit wide (LSB of the 24 on GDB) */

wire REPEAT;				/* REP instruction signal - generated by PCU */

wire AGU_C;					/* AGU generated carry bit that goes to the data ALU */

wire [7:0] CCR_from_alu;	/* condition code bits from the data alu */

wire [7:0] CCR;				/* the CCR register from the PCU */

wire Swrite;				/* S bit (in the CCR) write enable from the data alu */

wire Lwrite;				/* L bit (in the CCR) write enable from the data alu */

wor J;						/* jump bit that comes from either the AGU or the data ALU and goes to the PCU */


/*==============================================================================*/

/*===========	Module Instantiation	========================================*/

/*--------------------------*/
/*			AGU				*/
/*--------------------------*/

agu agu (
	.reset (reset),
	.PDB (PDB),
	.GDB (GDB),
	.REPEAT (REPEAT),
	.E (CCR[5]),
	.U (CCR[4]),
	.Z (CCR[2]),
	.PAB (PAB),
	.XAB (XAB),
	.YAB (YAB),
	.XWRITE (XWRITE),
	.XREAD  (XREAD),
	.YWRITE (YWRITE),
	.YREAD  (YREAD),
	.C (AGU_C),
	.J (J),
	.Clk (Clk)
	);


/*--------------------------*/
/*		data_alu			*/
/*--------------------------*/

data_alu data_alu (
	.reset (reset),
	.PDB (PDB),
	.XDB (XDB),
	.YDB (YDB),
	.REPEAT (REPEAT),
	.AGU_C (AGU_C),
	.S1 (S1),
	.S0 (S0),
	.CCR (CCR),
	.CCR_from_alu (CCR_from_alu),
	.Swrite (Swrite),
	.Lwrite (Lwrite),
	.J (J),
	.Clk (Clk)
	);


/*--------------------------*/
/*		bus_switch			*/
/*--------------------------*/

bus_switch bus_switch (
	.reset (reset),
	.PDB (PDB),
	.GDB (GDB),
	.XDB (XDB),
	.YDB (YDB),
	.REPEAT (REPEAT),
	.Clk (Clk)
	);


/*--------------------------*/
/*			PCU				*/
/*--------------------------*/

pcu PCU(
	.reset (reset),
	.PDB (PDB),
	.GDB (GDB_PCU),
	.PAB_in (PAB),
	.CCR_from_alu (CCR_from_alu),
	.Swrite (Swrite),
	.Lwrite (Lwrite),
	.J (J),
	.PAB_out (PAB),
	.REPEAT (REPEAT),
	.CCR (CCR),
	.S1 (S1),
	.S0 (S0),
	.Clk (Clk)
	);


/*==================================================*/


assign GDB_PCU = GDB[`addrbus];		/* the PCU loads only the 16-LSB of the GDB bus */




endmodule	/* core */
