/*	File:	shift1.v	  						*/

/*	module name: shift1						*/

/*	Description: 1 bit shifter module for ALU 		*/

/*				arithmatical shift one bit left or right		*/


/*==============================================================================*/


/********************************************************************************/
/*																				*/
/*	module:																		*/
/*																				*/
/********************************************************************************/

module shift1 (
	left, right,
	in,    /* in2, ext:msb:lsb */
	out
	);


/*============	I/O direction	================================================*/

input		left, right;
input [`acc]	in;
output [`acc]	out;

/*==============================================================================*/



/*============		I/O type	========================================*/

reg [`acc] out;		

/*==============================================================================*/


/*==============================================================================*/
/*	processes																	*/
/*==============================================================================*/


always @(left or right or in )
begin
	if (left)
		out = {in[54:0], 1'b0};
	else if (right)
		out = {in[55], in[55:1]};
	else
		out = in;
end   /* always */


endmodule	/* end module */
