/*	File:	core_test.v	  		*/

/*	module name: top				*/

/*	Description: TEST FILE			*/

/*	Tested Module name:	core.v		*/

/*	Author: Nitzan Weinberg */


/*==============================================================================*/

/********************************************************************************/
/*																				*/
/*	module:	top																	*/
/*																				*/
/********************************************************************************/

module top;



/*============		I/O type	================================================*/

reg reset;

reg [`databus] PDB;
wire [`databus] XDB;
wire [`databus] YDB;

wire [`addrbus] PAB;

wire [`addrbus] XAB;
wire Xwrite;
wire Xread;

wire [`addrbus] YAB;
wire Ywrite;
wire Yread;

reg Clk;


/*==============================================================================*/

/*============		 internal nets			=========*/

reg [`databus] XDB_in;
reg [`databus] YDB_in;




/*===========	Module Instantiations	 =======================================*/

core core(
	.reset  (reset),
	.PDB    (PDB),
	.XDB    (XDB),
	.YDB    (YDB),
	.PAB    (PAB),
	.XAB    (XAB),
	.XWRITE (XWRITE),
	.XREAD  (XREAD),
	.YAB    (YAB),
	.YWRITE (YWRITE),
	.YREAD  (YREAD),
	.Clk    (Clk)
	);


/*==============================================================================*/

/* XDB and YDB driven by the memories */

assign XDB = XDB_in;	/* driven by the X data memory */
assign YDB = YDB_in;	/* driven by the Y data memory */


/*==============================================================================*/
/*	initialize																		*/
/*==============================================================================*/

initial
	begin
		$shm_open("waves.shm");		/* generates a dump file for cWaves to use */

		$shm_probe("AS");			/* keep track of all signals in the current and lower modules in the hierarcy */
		
		
		Clk = 0;
		XDB_in = 24'hzzzzzz;
		YDB_in = 24'hzzzzzz;
		reset = 1;	/* for one clock cycle */
		
		#10 reset = 0;
		
		/* I: */

		    PDB = 24'b001_10_000_00000111_00000000; /* r0 = 7 */
		#10 PDB = 24'b001_10_110_00001111_00000000; /* r6 = f */
		#10 PDB = 24'b001_11_011_00011111_00000000; /* n3 = 1f */
		#10 PDB = 24'b001_11_110_00111111_00000000; /* n6 = 3f */

		/* 40 */

		/* R: */

		/* from agu to data alu */
		
		#10 PDB = 24'b001000_10_000_00_100_00000000; /* r0 -> x0 = 7 */
		
		#10 PDB = 24'b001000_10_110_00_111_00000000; /* r6 -> y1 = f */

		#10 PDB = 24'b001000_11_011_01_001_00000000; /* n3 -> b0 = 1f */

		#10 PDB = 24'b001000_11_110_01_010_00000000; /* n6 -> a2 = 3f */

		/* 80 */
		
		/* from agu to agu */
		
		#10 PDB = 24'b001000_10_000_10_001_00000000; /* r0 -> r1 = 7 */

		#10 PDB = 24'b001000_10_110_10_011_00000000; /* r6 -> r3 = f */
		
		#10 PDB = 24'b001000_10_001_11_010_00000000; /* r1 -> n2 = 7 */

		#10 PDB = 24'b001000_10_011_11_111_00000000; /* r3 -> n7 = f */

		#10 PDB = 24'b001000_11_011_11_001_00000000; /* n3 -> n1 = 1f */

		#10 PDB = 24'b001000_11_110_10_111_00000000; /* r6 -> r7 = 3f */

		#10 PDB = 24'b001000_11_010_10_010_00000000; /* n2 -> r2 = 7 */

		#10 PDB = 24'b001000_11_111_10_100_00000000; /* n7 -> r4 = f */

		#10 PDB = 24'b001000_11_001_10_101_00000000; /* n1 -> r5 = 1f */

		/* 170 */
		
		/* from data alu to data alu */
		
		#10 PDB = 24'b001000_00_100_00_101_00000000; /* x0 -> x1 = 7 */

		#10 PDB = 24'b001000_00_101_00_110_00000000; /* x1 -> y0 = 7 */
		
		#10 PDB = 24'b001000_00_100_01_101_00000000; /* x0 -> b1 = 7 */

		#10 PDB = 24'b001000_00_110_01_100_00000000; /* y0 -> a1 = 7 */

		#10 PDB = 24'b001000_00_111_01_011_00000000; /* y1 -> b2 = f */

		#10 PDB = 24'b001000_01_001_01_000_00000000; /* b0 -> a0 = 1f */


		#10 PDB = 24'b001000_01_000_00_100_00000000; /* a0 -> x0 = 1f */
		
		#10 PDB = 24'b001000_01_100_00_111_00000000; /* a1 -> y1 = 7 */

		#10 PDB = 24'b001000_01_010_01_100_00000000; /* a2 -> a1 = 3f */

		#10 PDB = 24'b001000_01_001_00_110_00000000; /* b0 -> y0 = 1f */

		#10 PDB = 24'b001000_00_110_00_111_00000000; /* y0 -> y1 = 1f */

		/* 280 */
		
		/* data alu to agu */
		
		#10 PDB = 24'b001000_00_100_10_001_00000000; /* x0 -> r1 = 1f */

		#10 PDB = 24'b001000_01_010_11_101_00000000; /* a2 -> n5 = 3f */

		#10 PDB = 24'b001000_00_111_10_011_00000000; /* y1 -> r3 = 1f */

		#10 PDB = 24'b001000_01_101_10_100_00000000; /* b1 -> r4 = 7 */

		/* 320 */
		
		/* agu to data alu */

		#10 PDB = 24'b001000_11_101_00_101_00000000; /* n5 -> x1 = 3f */

		#10 PDB = 24'b001000_11_010_01_001_00000000; /* n2 -> b0 = 7 */

		#10 PDB = 24'b001000_10_111_00_111_00000000; /* r7 -> y1 = 3f */

		#10 PDB = 24'b001000_10_001_01_010_00000000; /* r1 -> a2 = 1f */

		/* 360 */
		
		/* U: */

		/*                        MM RRR              */
		#10 PDB = 24'b00100000010_00_011_00000000; /* (r3)-n3 -> r3 = 0 */

		#10 PDB = 24'b00100000010_11_011_00000000; /* (r3)+ -> r3 = 1 */

		#10 PDB = 24'b00100000010_01_010_00000000; /* (r2)+n2 -> r2 = e */

		#10 PDB = 24'b00100000010_10_010_00000000; /* (r2)- -> r2 = d */

		#10 PDB = 24'b00100000010_11_110_00000000; /* (r6)+ -> r6 = 10 */

		#10 PDB = 24'b00100000010_10_100_00000000; /* (r4)- -> r4 =  6 */

		
		/* 420 */
		
		
		/* X: or Y: */

		/* type I */
		/*					X							*/
		/*               dd Y ddd W F MMM RRR			*/  
		#10 PDB = 24'b01_00_0_100_1_1_000_010_00000000; /* x:(r2)-n2, x0 */

		#10 PDB = 24'b01_11_1_100_1_1_011_111_00000000; /* y:(r7)+, n4 */
		    
		#10	PDB = 24'h000000;
			XDB_in = 24'h100;

		#10 PDB = 24'b01_00_0_111_1_1_101_100_00000000; /* x:(r4+n4), y1 */
			YDB_in = 24'h200;
			XDB_in = 24'hzzzzzz;
			
		#10	PDB = 24'b01_00_0_100_0_1_011_011_00000000; /* x0, x:(r3)+ */
			YDB_in = 24'hzzzzzz;
		    
		#10 PDB = 24'b01_10_0_010_0_1_111_010_00000000; /* r2, x:-(r2) */
			XDB_in = 24'h300;

		/* type II */

		#10 PDB = 24'b01_00_1_101_1_0_000100_00000000;  /* y:4, x1 */
			XDB_in = 24'hzzzzzz;

		#10 PDB = 24'b01_10_1_101_0_0_000111_00000000;  /* r5, y:7 */
		
		#10	PDB = 24'h000000;
			YDB_in = 24'h400;


		/* 510 */
		
		/* X:R Class I */

		/*                 ff d f W   MMM RRR			*/  
		#10 PDB = 24'b0001_00_1_1_0_0_001_111_00000000; /* x0, x:(r7)+n7  B -> y1 */
			YDB_in = 24'hzzzzzz;
		
		#10 PDB = 24'b0001_10_1_0_0_0_011_010_00000000; /* A, x:(r2)+  B -> y0 */

		
		/* 530ns */
		

		/* X:Y: */
		
		/*              w mm ee ff W rr MM RRR          */
		#10 PDB = 24'b1_1_10_01_01_0_11_11_111_00000000; /* x1, x:(r7)+  y:(r3)-, y1*/

		#10 PDB = 24'h000000;
		
		#10	YDB_in = 24'h2000;

		/* 560 */


		/* X: or Y: */

		/* immediate data */

		/*					X						*/
		/*               dd Y ddd W F MMM RRR			*/  

		#10 PDB = 24'b01_11_1_000_1_1_110_100_00000000; /* y:imm, n0 */
			YDB_in = 24'hzzzzzz;
		
		#10 PDB = 24'h500;

		#10 PDB = 24'b01_11_1_101_0_1_001_011_00000000; /* n5, y:(r3)+n3 */

		#10 PDB = 24'b01_11_0_000_0_1_010_100_00000000; /* n0, x:(r4)- */


		/* 600ns */


		/* X: or Y: */
		
		/* absolute address */

		/*					X						*/
		/*               dd Y ddd W F MMM RRR			*/  

		#10 PDB = 24'b01_11_1_110_1_1_110_000_00000000; /* y:abs, n6 */
		
		#10 PDB = 24'h44;

		#10	YDB_in = 24'hB; PDB = 24'h000000;

		#10	YDB_in = 24'hzzzzzz;
			


		/* R:Y Class I */
		
		/* immediate data */
		
		
		/*                 d e ff W   MMM RRR			*/  
		#10	PDB = 24'b0001_0_0_00_1_1_110_100_00000000; /* A:x0  imm,y0 */
					
		#10 PDB = 24'hA;
		
		/* 640ns */


		#10 PDB = 24'h000000;

/*============================================================*/
		

		/* immediate data X: type 1 */

		/*					X						*/
		/*               dd Y ddd W F MMM RRR			*/  

//		#10 PDB = 24'b01_00_0_100_1_1_110_100_00000000; /* x0 */
		
//		#10 PDB = 24'h123456;

//		#10 PDB = 24'b01_00_0_101_1_1_110_100_00000000; /* x1 */
		
//		#10 PDB = 24'h3;

//		#10 PDB = 24'b01_00_0_110_1_1_110_100_00000000; /* y0 */
		
//		#10 PDB = 24'h654321;

//		#10 PDB = 24'b01_00_0_111_1_1_110_100_00000000; /* y1 */
		
//		#10 PDB = 24'h654321;

//		#10 PDB = 24'b01_01_0_100_1_1_110_100_00000000; /* a1 */
		
//		#10 PDB = 24'h020304;

//		#10 PDB = 24'b01_01_0_000_1_1_110_100_00000000; /* a0 */
		
//		#10 PDB = 24'h0;

//		#10 PDB = 24'b01_01_0_101_1_1_110_100_00000000; /* b1 */
		
//		#10 PDB = 24'h123456;

//		#10 PDB = 24'b01_01_0_001_1_1_110_100_00000000; /* b0 */
		
//		#10 PDB = 24'h789abc;


		/* 760ns */
		
		
		/* I */
		#10 PDB = 24'b001_01010_00000000_00000000; /* a2 */
		#10 PDB = 24'b001_01100_00000000_00000000; /* a1 */
		#10 PDB = 24'b001_01000_00000001_00000000; /* a0 */

//		#10 PDB = 24'b001_01011_00000000_00000000; /* b2 */
//		#10 PDB = 24'b001_01101_10000000_00000000; /* b1 */
//		#10 PDB = 24'b001_01001_00000001_00000000; /* b0 */
		
//		#10 PDB = 24'b001_10011_00000000_00000000; /* R3 */



		/* I */

//		#10 PDB = 24'b001_10010_01001011_00000000; /* R2 = 4B */

//		#10 PDB = 24'b001_11100_00000110_00000000; /* n4 = 6 */
		

		/* U: */
		/*                        MM RRR              */
//		#10 PDB = 24'b00100000010_01_100_00000000; /* (r4)+n4 */


		/* L: */
		/*                 L   LL W F MMMRRR         */
//		#10 PDB = 24'b0100_0_0_10_0_1_011000_00000000;	/* X, L:(r0)+ */

//		#10 PDB = 24'b0100_0_0_01_1_1_010000_00000000;	/* L:(r0)-, B10 */

//		#10 PDB = 24'h000000;
		
//		#10 XDB_in = 24'h111; YDB_in = 24'hfff222;
		
//		#10 XDB_in = 24'hzzzzzz; YDB_in = 24'hzzzzzz;
		
			/* absolute address */
//		#10 PDB = 24'b0100_1_0_11_0_1_011000_00000000;	/* BA, L:(r0)+ */

//		#10 PDB = 24'b0100_1_0_00_1_1_110000_00000000;	/* L:75, A */

//		#10 PDB = 24'h75;	/* absolute addr */
		
//		#10 XDB_in = 24'hfff333; YDB_in = 24'h444;
//			PDB = 24'h000000;
		
//		#10 XDB_in = 24'hzzzzzz; YDB_in = 24'hzzzzzz;



		/* I */

//		#10 PDB = 24'b001_10010_01001011_00000000; /* R2 = 4B */

//		#10 PDB = 24'b001_11010_00000010_00000000; /* n2 = 2 */

//		#10 PDB = 24'b001_10100_00000101_00000000; /* R4 = 5 */

//		#10 PDB = 24'b001_11100_00000011_00000000; /* n4 = 3 */

//		#10 PDB = 24'b001_10111_11111111_00000000; /* R7 = FF */

//		#10 PDB = 24'b001_11111_11111111_00000000; /* n7 = FF */



		#10 PDB = 24'h000000;
		#10 PDB = 24'h000000;
		

		/* LUA */
		/*                         MM RRR      dddd  */
//		#10 PDB = 24'b00000100_010_11_010_0001_0011;	/* LUA (r0)+n0 -> r1 */




`ifdef test
		/* DO Class III */
		/*                     iiiiiiii      hhhh  */
		#10 PDB = 24'b00000110_00000011_1000_0000;	/* DO #3, expr */
		
		#10 PDB = 24'h4c;	/* expr (first inst address after the end of the loop) */

		
		/* U: */
		/*                        MM RRR              */
		#10 PDB = 24'b00100000010_01_010_00000000; /* (r2)+n2 */

		#10 PDB = 24'b00100000010_01_100_00000000; /* (r4)+n4 */

		#10 PDB = 24'b00100000010_01_111_00000000; /* (r7)+n7 */

		#10 PDB = 24'b00100000010_01_010_00000000; /* (r2)+n2 */

		#10 PDB = 24'b00100000010_01_100_00000000; /* (r4)+n4 */

		#10 PDB = 24'b00100000010_01_111_00000000; /* (r7)+n7 */

		#10 PDB = 24'b00100000010_01_010_00000000; /* (r2)+n2 */

		#10 PDB = 24'b00100000010_01_100_00000000; /* (r4)+n4 */

		#10 PDB = 24'b00100000010_01_111_00000000; /* (r7)+n7 */

		#10 PDB = 24'b00100000010_01_010_00000000; /* (r2)+n2 */

		#10 PDB = 24'b00100000010_01_100_00000000; /* (r4)+n4 */

		#10 PDB = 24'b00100000010_01_111_00000000; /* (r7)+n7 */
`endif



`ifdef test
		/* DO Class IV */
		/*                        DDDDDD     	  */
		#10 PDB = 24'b00000110_11_100101_00000000;	/* DO m5, expr */
		
		#10 PDB = 24'h4d;	/* expr (first inst address after the end of the loop) */

		
		/* U: */
		/*                        MM RRR              */
		#10 PDB = 24'b00100000010_01_010_00000000; /* (r2)+n2 */

		#10 PDB = 24'b00100000010_01_100_00000000; /* (r4)+n4 */

		#10 PDB = 24'b00100000010_01_111_00000000; /* (r7)+n7 */

		#10 PDB = 24'b00100000010_01_010_00000000; /* (r2)+n2 */

		#10 PDB = 24'b00100000010_01_100_00000000; /* (r4)+n4 */

		#10 PDB = 24'b00100000010_01_111_00000000; /* (r7)+n7 */

		#10 PDB = 24'b00100000010_01_010_00000000; /* (r2)+n2 */

		#10 PDB = 24'b00100000010_01_100_00000000; /* (r4)+n4 */

		#10 PDB = 24'b00100000010_01_111_00000000; /* (r7)+n7 */

		#10 PDB = 24'b00100000010_01_010_00000000; /* (r2)+n2 */

		#10 PDB = 24'b00100000010_01_100_00000000; /* (r4)+n4 */

		#10 PDB = 24'b00100000010_01_111_00000000; /* (r7)+n7 */

		#10 PDB = 24'b00100000010_01_010_00000000; /* (r2)+n2 */

		#10 PDB = 24'b00100000010_01_100_00000000; /* (r4)+n4 */

		#10 PDB = 24'b00100000010_01_111_00000000; /* (r7)+n7 */

		#10 PDB = 24'b00100000010_01_010_00000000; /* (r2)+n2 */

		#10 PDB = 24'b00100000010_01_100_00000000; /* (r4)+n4 */

		#10 PDB = 24'b00100000010_01_111_00000000; /* (r7)+n7 */

		#10 PDB = 24'b00100000010_01_010_00000000; /* (r2)+n2 */

		#10 PDB = 24'b00100000010_01_100_00000000; /* (r4)+n4 */

		#10 PDB = 24'b00100000010_01_111_00000000; /* (r7)+n7 */
`endif






		/* X: or Y: */

		/* type I */
		/*					X							*/
		/*               dd Y ddd W F MMM RRR			*/  
//		#10 PDB = 24'b01_11_0_001_0_1_001_000_00000000; /* n1, x:(r0)+n0 */



// ***********************************************
// testing nested loops for sphinx3 
// ***********************************************
`ifdef test
		/* I */
		/*                ddddd iiiiiiii			*/
		#10 PDB = 24'b001_10000_00000000_00000000; /* r0 = 0 */

		#10 PDB = 24'b001_11000_00010000_00000000; /* n0 = 10 */

		#10 PDB = 24'b001_10001_00000000_00000000; /* r1 = 0 */

		#10 PDB = 24'b001_11001_00010000_00000000; /* n1 = 10 */

		#10 PDB = 24'b001_10111_00000000_00000000; /* r7 = 0 */

		#10 PDB = 24'b001_11111_00010000_00000000; /* n7 = 10 */

		#10 PDB = 24'b001_10101_00000000_00000000; /* r5 = 0 */

		#10 PDB = 24'b001_11101_00010000_00000000; /* n5 = 10 */

		#10 PDB = 24'b001_10110_00000000_00000000; /* r6 = 0 */

		#10 PDB = 24'b001_11110_00010000_00000000; /* n6 = 10 */

		#10 PDB = 24'b001_10010_00000000_00000000; /* r2 = 0 */

		#10 PDB = 24'b001_11010_00010000_00000000; /* n2 = 10 */

		#10 PDB = 24'b001_10100_00000000_00000000; /* r4 = 0 */

		#10 PDB = 24'b001_10011_00000000_00000000; /* r3 = 0 */



		/* DO Class III */
		/*                     iiiiiiii      hhhh  */
		#10 PDB = 24'b00000110_00001000_1000_0000;	/* DO #8, expr    pc=55 */
		
		#10 PDB = 24'h63;	/* expr (first inst address after the end of the loop) */


		/* --- begin outer loop itteration 1 --- */
		
		/* X:Y: */
		/*              w mm ee ff W rr MM RRR          */
		#10 PDB = 24'b1_1_11_01_10_1_00_11_000_00000000; /* x:(r0)+,x1  y:(r4)+, A   pc=57*/



		/* DO Class III */
		/*                     iiiiiiii      hhhh  */
		#10 PDB = 24'b00000110_00000011_1000_0000;	/* DO #3, expr   pc=58 */
		
		#10 PDB = 24'h62;	/* expr (first inst address after the end of the loop) */


		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 1 - pc=61*/

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 2 - pc=61 */

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 3 - pc=61 */

		#10 PDB = 24'h000001;   /* end of outer loop - itteration 1 - pc=62 */


		/* --- begin outer loop itteration 2 --- */

		
		/* X:Y: */
		/*              w mm ee ff W rr MM RRR          */
		#10 PDB = 24'b1_1_11_01_10_1_00_11_000_00000000; /* x:(r0)+,x1  y:(r4)+, A   pc=57*/



		/* DO Class III */
		/*                     iiiiiiii      hhhh  */
		#10 PDB = 24'b00000110_00000011_1000_0000;	/* DO #3, expr   pc=58 */
		
		#10 PDB = 24'h62;	/* expr (first inst address after the end of the loop) */


		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 1 - pc=61*/

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 2 - pc=61 */

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 3 - pc=61 */

		#10 PDB = 24'h000001;   /* end of outer loop - itteration 2 - pc=62 */


		/* --- begin outer loop itteration 3 --- */

		
		/* X:Y: */
		/*              w mm ee ff W rr MM RRR          */
		#10 PDB = 24'b1_1_11_01_10_1_00_11_000_00000000; /* x:(r0)+,x1  y:(r4)+, A   pc=57*/



		/* DO Class III */
		/*                     iiiiiiii      hhhh  */
		#10 PDB = 24'b00000110_00000011_1000_0000;	/* DO #3, expr   pc=58 */
		
		#10 PDB = 24'h62;	/* expr (first inst address after the end of the loop) */


		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 1 - pc=61*/

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 2 - pc=61 */

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 3 - pc=61 */

		#10 PDB = 24'h000001;   /* end of outer loop - itteration 3 - pc=62 */


		/* --- begin outer loop itteration 4 --- */

		
		/* X:Y: */
		/*              w mm ee ff W rr MM RRR          */
		#10 PDB = 24'b1_1_11_01_10_1_00_11_000_00000000; /* x:(r0)+,x1  y:(r4)+, A   pc=57*/



		/* DO Class III */
		/*                     iiiiiiii      hhhh  */
		#10 PDB = 24'b00000110_00000011_1000_0000;	/* DO #3, expr   pc=58 */
		
		#10 PDB = 24'h62;	/* expr (first inst address after the end of the loop) */


		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 1 - pc=61*/

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 2 - pc=61 */

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 3 - pc=61 */

		#10 PDB = 24'h000001;   /* end of outer loop - itteration 3 - pc=62 */


		/* --- begin outer loop itteration 5 --- */

		
		/* X:Y: */
		/*              w mm ee ff W rr MM RRR          */
		#10 PDB = 24'b1_1_11_01_10_1_00_11_000_00000000; /* x:(r0)+,x1  y:(r4)+, A   pc=57*/



		/* DO Class III */
		/*                     iiiiiiii      hhhh  */
		#10 PDB = 24'b00000110_00000011_1000_0000;	/* DO #3, expr   pc=58 */
		
		#10 PDB = 24'h62;	/* expr (first inst address after the end of the loop) */


		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 1 - pc=61*/

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 2 - pc=61 */

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 3 - pc=61 */

		#10 PDB = 24'h000001;   /* end of outer loop - itteration 3 - pc=62 */


		/* --- begin outer loop itteration 6 --- */

		
		/* X:Y: */
		/*              w mm ee ff W rr MM RRR          */
		#10 PDB = 24'b1_1_11_01_10_1_00_11_000_00000000; /* x:(r0)+,x1  y:(r4)+, A   pc=57*/



		/* DO Class III */
		/*                     iiiiiiii      hhhh  */
		#10 PDB = 24'b00000110_00000011_1000_0000;	/* DO #3, expr   pc=58 */
		
		#10 PDB = 24'h62;	/* expr (first inst address after the end of the loop) */


		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 1 - pc=61*/

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 2 - pc=61 */

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 3 - pc=61 */

		#10 PDB = 24'h000001;   /* end of outer loop - itteration 3 - pc=62 */


		/* --- begin outer loop itteration 7 --- */

		
		/* X:Y: */
		/*              w mm ee ff W rr MM RRR          */
		#10 PDB = 24'b1_1_11_01_10_1_00_11_000_00000000; /* x:(r0)+,x1  y:(r4)+, A   pc=57*/



		/* DO Class III */
		/*                     iiiiiiii      hhhh  */
		#10 PDB = 24'b00000110_00000011_1000_0000;	/* DO #3, expr   pc=58 */
		
		#10 PDB = 24'h62;	/* expr (first inst address after the end of the loop) */


		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 1 - pc=61*/

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 2 - pc=61 */

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 3 - pc=61 */

		#10 PDB = 24'h000001;   /* end of outer loop - itteration 3 - pc=62 */


		/* --- begin outer loop itteration 8 --- */

		
		/* X:Y: */
		/*              w mm ee ff W rr MM RRR          */
		#10 PDB = 24'b1_1_11_01_10_1_00_11_000_00000000; /* x:(r0)+,x1  y:(r4)+, A   pc=57*/



		/* DO Class III */
		/*                     iiiiiiii      hhhh  */
		#10 PDB = 24'b00000110_00000011_1000_0000;	/* DO #3, expr   pc=58 */
		
		#10 PDB = 24'h62;	/* expr (first inst address after the end of the loop) */


		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 1 - pc=61*/

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 2 - pc=61 */

		#10 PDB = 24'h21cf00;
		
		#10 PDB = 24'hf5b964;
		
		#10 PDB = 24'h11de7c;

		#10 PDB = 24'h21e680;
		
		#10 PDB = 24'h12e798;
		
		#10 PDB = 24'h1ea2a2;
		
		#10 PDB = 24'h86f8ba;

		#10 PDB = 24'hfe0200;	/* end inner loop - itteration 3 - pc=61 */

		#10 PDB = 24'h000001;   /* end of outer loop - itteration 3 - pc=62 */



		#10 PDB = 24'h000010;	/* sp=63 */

		#10 PDB = 24'h000100;	/* sp=64 */

		#10 PDB = 24'h001000;	/* sp=65 */
`endif

// ***********************************************

		/* ABS */
		/*                                   d       */
//		#10 PDB = 24'b00000000_00000000_0010_0_110;


		/* ADD */
//		#10 PDB = 24'b00000000_00000000_0_100_0_000;


		/* ADDL */
		/*                                   d       */
//		#10 PDB = 24'b00000000_00000000_0001_1_010;


		/* AND */
		/*                                 JJ d       */
//		#10 PDB = 24'b00000000_00000000_01_00_0_110;


		/* ANDI */
		/*                     iiiiiiii        EE    */
//		#10 PDB = 24'b00000000_11111100_101110_10;


		/* ASL */
		/*                                   d       */
//		#10 PDB = 24'b00000000_00000000_0011_0_010;


		/* ASR */
		/*                                   d       */
//		#10 PDB = 24'b00000000_00000000_0010_1_010;


		/*---------*/
		/* B C L R */
		/*---------*/

		/* BCLR I */
		/*                        MMM RRR   S   bbbbb   */
//		#10 PDB = 24'b00001010_01_101_110_0_1_0_00101; /* #5, y:(r6+n6) */
		
//		#10 PDB = 24'h000000;

//		#10	YDB_in = 24'h888828;	/* will change to 888808 */

//		#10	YDB_in = 24'hzzzzzz;

			/* absolute address */
//		#10 PDB = 24'b00001010_01_110_000_0_1_0_00101; /* #5, y:#2323 */
		
//		#10 PDB = 24'hbb2323;	/* addr */

//		#10	YDB_in = 24'h888828;	/* will change to 888808 */
//			PDB = 24'h000000;

//		#10	YDB_in = 24'hzzzzzz;
		

		/* BCLR II */
		/*                        aaaaaa   S   bbbbb   */
//		#10	PDB = 24'b00001010_00_000100_0_0_0_00000; /* #0, x:4 */

//		#10 PDB = 24'h000000;

//		#10	XDB_in = 24'ha44447;	/* will change to a44446 */

//		#10	XDB_in = 24'hzzzzzz;


		/* BCLR III */
		/*                        DDD_DDD     bbbbb   */
//		#10	PDB = 24'b00001010_11_010_000_010_00000;	/* r0 = 6 */

//		#10 PDB = 24'b00001010_11_011_010_010_00010;	/* n2 = 3 */

//		#10 PDB = 24'h000000;
		
//		#10 PDB = 24'b01_11_0_111_0_1_101_010_00000000;	/* move n7->X:(r2+n2)*/
		
//		#10 PDB = 24'b00001010_11_001_000_010_00001;	/* a0 = 1D */

//		#10 PDB = 24'b00001010_11_001_011_010_00001;	/* b2 = D */

//		#10 PDB = 24'b00001010_11_000_111_010_00000;	/* y1 = 2000 */

//		#10 PDB = 24'b00001010_11_111_001_010_01001;	/* I1 = 0 */

//		#10 PDB = 24'b00001010_11_001_111_010_00111;	/* B = _ff7f */

//		#10 PDB = 24'b00001010_11_001_111_010_00110;	/* B = no effect */



		/*---------*/
		/* B S E T */
		/*---------*/

		/* BSET I */
		/*                        MMM RRR   S   bbbbb   */
//		#10 PDB = 24'b00001010_01_101_110_0_1_1_00101;	/* #5, y:(r6+n6) */
		
//		#10 PDB = 24'h000000;
		
//		#10	YDB_in = 24'h888888; /* will change to 8888A8 */

//			PDB = 24'b00001010_01_110_000_0_1_1_01000;	/* y:abs addr */

//		#10	YDB_in = 24'hzzzzzz;

//			PDB = 24'heee;

//		#10 YDB_in = 24'he00; /* will change to F00 */
//			PDB = 24'h000000;	/* no need for this if next inst is used */

//		#10 YDB_in = 24'hzzzzzz;


		/* BSET II */
		/*                        aaaaaa   S   bbbbb   */
//			PDB = 24'b00001010_00_001000_0_0_1_00000; /* #0, x:$8 */

//		#10 PDB = 24'h000000;

//		#10	XDB_in = 24'ha44446; /* will change to A44447 */

//		#10	XDB_in = 24'hzzzzzz;

		/* BSET III */
		/*                        DDD_DDD     bbbbb   */
//			PDB = 24'b00001010_11_010_000_011_00100;	/* r0 = 17 */

//		#10 PDB = 24'b00001010_11_011_010_011_00010;	/* n2 = 7 no change */

//		#10 PDB = 24'h000000;
		
//		#10 PDB = 24'b01_11_0_111_0_1_101_010_00000000;	/* move n7->X:(r2+n2)*/
		
//		#10 PDB = 24'b00001010_11_001_000_011_00101;	/* a0 = 3F */

//		#10 PDB = 24'b00001010_11_001_011_011_00100;	/* b2 = 1F */

//		#10 PDB = 24'b00001010_11_000_111_011_00000;	/* y1 = 2001 */

//		#10 PDB = 24'b00001010_11_111_001_011_01001;	/* I1 = 1 no change */

//		#10 PDB = 24'b00001010_11_001_111_011_00111;	/* B = 7fffff */

//		#10 PDB = 24'b00001010_11_001_111_011_00110;	/* B no effect */

//		#10 PDB = 24'b00001010_11_000_101_011_10111;	/* x1 800400 */


		/*---------*/
		/* B T S T */
		/*---------*/

		/* BTST I */
		/*                        MMM RRR   S   bbbbb   */
//		#10 PDB = 24'b00001011_01_101_110_0_1_1_00101;	/* #5, y:(r6+n6) */
		
//		#10 PDB = 24'h000000;

//		#10	YDB_in = 24'h8888a8; /* C = 1 */
//			PDB = 24'b00001011_01_110_000_0_1_1_01000;	/* #8, y:abs addr */

//		#10 PDB = 24'heee;
//			YDB_in = 24'hzzzzzz;

//		#10 YDB_in = 24'hf00; /* C = 1 */
//			PDB = 24'h000000;

		/* BTST II */
		/*                        aaaaaa   S   bbbbb   */
//		#10	PDB = 24'b00001011_00_001000_0_0_1_00000; /* #0, x:$8 */
//			YDB_in = 24'hzzzzzz;

//		#10 PDB = 24'h000000;

//		#10	XDB_in = 24'ha44447; /* C = 1 */
		
//		#10 XDB_in = 24'hzzzzzz;


		/* BTST III */
		/*                        DDD_DDD     bbbbb   */
//			PDB = 24'b00001011_11_010_000_011_00000;	/* r0, C = 1 */

//		#10 PDB = 24'b00001011_11_011_010_011_00010;	/* n2, C = 1 */

//		#10 PDB = 24'h000000;
		
//		#10 PDB = 24'b01_11_0_111_0_1_101_010_00000000;	/* move n7->X:(r2+n2)*/
		
//		#10 PDB = 24'b00001011_11_001_000_011_00001;	/* a0, C = 1 */

//		#10 PDB = 24'b00001011_11_001_011_011_00001;	/* b2, C = 1 */

//		#10 PDB = 24'b00001011_11_000_111_011_00000;	/* y1, C = 0 */

//		#10 PDB = 24'b00001011_11_111_001_011_01001;	/* I1, C = 1 */

//		#10 PDB = 24'b00001011_11_001_111_011_00111;	/* B=7fffff, C = 1 */

//		#10 PDB = 24'b00001011_11_001_111_011_00110;	/* B no effect */

//		#10 PDB = 24'b00001011_11_000_101_011_10111;	/* x1, C = 0 */


		/* CLR */
		/*                                   d       */
//		#10 PDB = 24'b00000000_00000000_0001_0_011;


		/* CMP */
		/*                       JJJ d               */
//		#10 PDB = 24'b00000000_0_101_1_101;


		/* CMPM */
		/*                       JJJ d               */
//		#10 PDB = 24'b00000000_0_110_0_111;


		/* EOR */
		/*                                 JJ d       */
//		#10 PDB = 24'b00000000_00000000_01_11_1_011;


		/*---------*/
		/* J C L R */
		/*---------*/

		/* JCLR Class I */
		/*                        MMM RRR   S   bbbbb     */
//		#10 PDB = 24'b00001010_01_011_000_1_0_0_00010; /* #2, x:(r0)+ */
//		#10 PDB = 24'h001111; /* abs addr to jump to */

//		#10 XDB_in = 24'h83; /* J = 0 */
//			PDB = 24'h000000;

//		#10 XDB_in = 24'hzzzzzz;


		/* JCLR Class II */
		/*                        aaaaaa   S   bbbbb     */
//			PDB = 24'b00001010_00_100000_1_1_0_10111; /* #23, y:$20 */
//		#10 PDB = 24'h002222; /* abs addr to jump to */

//		#10 YDB_in = 24'h700000; /* J = 0 */
//			PDB = 24'h000000;
		
//		#10 YDB_in = 24'hzzzzzz;


		/* JCLR Class III */
		/*                        DDDDDD     bbbbb     */
//		#10	PDB = 24'b00001010_11_000110_000_10111;	/* #23, y0, J = 0 */
//		#10 PDB = 24'h003333; /* abs addr to jump to */

//		#10 PDB = 24'b00001010_11_001100_000_00001;	/* #1, a1, J = 1 */
//		#10 PDB = 24'h004444; /* abs addr to jump to */

//		#10 PDB = 24'b00001010_11_010101_000_00110;	/* #6, r5, J = 0 */
//		#10 PDB = 24'h005555; /* abs addr to jump to */



		/* JMP Class I */
		/*                          aaaa aaaaaaaa   */
`ifdef test
		#10 PDB = 24'b00001100_0000_0000_00000110;

		#10 PDB = 24'h111111;
		
		#10 PDB = 24'h222222;

		#10 PDB = 24'h333333;
`endif



		/* JMP Class II */
		/*                        MMM RRR            */
			/* absolute */
`ifdef test
		#10 PDB = 24'b00001010_11_110_000_10000000;

		#10 PDB = 24'h010ccc; /* abs addr to jump to */

		#10 PDB = 24'h000111;

		#10 PDB = 24'b00001010_11_111_001_10000000;		/* jmp -(r1) */

		#10 PDB = 24'h001000;
		
		#10 PDB = 24'h002000;
`endif

		
		/*---------*/
		/* J S E T */
		/*---------*/
		
		/* JSET Class I */
		/*                        MMM RRR   S   bbbbb     */
`ifdef test
		#10 PDB = 24'b00001010_01_010_000_1_1_1_00010; /* #2, y:(r0)- */
		#10 PDB = 24'h006666; /* abs addr to jump to */

		#10	YDB_in = 24'hffc;	/* J = 1 */
			PDB = 24'h111000;

		#10	YDB_in = 24'hzzzzzz;
			PDB = 24'h222000;
`endif
			
			
		/* JSET Class II */
		/*                        aaaaaa   S   bbbbb     */
//		#10	PDB = 24'b00001010_00_110000_1_0_1_00000;
//		#10 PDB = 24'h007777;	/* abs addr to jump to */

//		#10 YDB_in = 24'hzzzzzz;
//		    XDB_in = 24'hc; 	/* J = 0 */
//		    PDB = 24'h000000;


		/* JSET Class III */
		/*                        DDDDDD     bbbbb     */
//		#10 PDB = 24'b00001010_11_000100_001_01010;	/* x0, J = 1 */
//			XDB_in = 24'hzzzzzz;
//		#10 PDB = 24'h008888; /* abs addr to jump to */

//		#10 PDB = 24'b00001010_11_001011_001_00000;	/* b2, J = 1 */
//		#10 PDB = 24'h009999; /* abs addr to jump to */

//		#10 PDB = 24'b00001010_11_011100_001_01111;	/* n4, J = 0 */
//		#10 PDB = 24'h00aaaa; /* abs addr to jump to */

//		#10 PDB = 24'b00001010_11_001110_001_10110;	/* A, J = 1 */
//		#10 PDB = 24'h00bbbb; /* abs addr to jump to */


		/* LSL */
		/*                                   d       */
//		#10 PDB = 24'b00000000_00000000_0011_1_011;


		/* LSR */
		/*                                   d       */
//		#10 PDB = 24'b00000000_00000000_0010_0_011;


		/* MAC Format 1 */
		/*                                QQQ d k     */
//		#10 PDB = 24'b00000000_00000000_1_000_0_0_10;


		/* MAC Format 2 */
		/*                         sssss    QQ d k     */
//		#10 PDB = 24'b00000001_000_00011_11_01_0_0_10;


		/* MACR Format 1 */
		/*                                QQQ d k     */
//		#10 PDB = 24'b00000000_00000000_1_101_1_0_11;


		/* MACR Format 2 */
		/*                         sssss    QQ d k     */
//		#10 PDB = 24'b00000001_000_01010_11_10_1_1_11;


		/* MPY Format 1 */
		/*                                QQQ d k     */
//		#10 PDB = 24'b00000000_00000000_1_111_0_1_00;


		/* MPY Format 2 */
		/*                         sssss    QQ d k     */
//		#10 PDB = 24'b00000001_000_01001_11_11_0_0_00;


		/* MPYR Format 1 */
		/*                                QQQ d k     */
//		#10 PDB = 24'b00000000_00000000_1_001_1_1_01;


		/* MPYR Format 2 */
		/*                         sssss    QQ d k     */
//		#10 PDB = 24'b00000001_000_01110_11_00_1_1_01;



		/* MOVEC Class I */
		/*                     W   MMMRRR   s   ddddd */
// 		#10 PDB = 24'b00000101_0_1_011001_0_0_1_00010;	/* m2, x:(r1)+ */

//		#10 PDB = 24'b00000101_1_1_101111_0_1_1_00010;	/* y:(r7+n7), m2 */

// 		#10 PDB = 24'h000000;
		
// 		#10 YDB_in = 24'h88aaaa;
		
// 		#10 PDB = 24'b00000101_0_1_111111_0_0_1_00010;	/* m2, x:-(r7) */
// 			YDB_in = 24'hzzzzzz;

// 		#10 PDB = 24'h000000;

			/* immediate data */
// 		#10 PDB = 24'b00000101_1_1_110100_0_0_1_00100;	/* #008003, m4 */

//		#10 PDB = 24'h008003;
		
// 		#10	PDB = 24'b00000101_0_1_011001_0_0_1_00100;	/* m4, x:(r1)+ */

			/* absolute address */
// 		#10 PDB = 24'b00000101_1_1_110000_0_1_1_00000;	/* y:#12, m0 */

// 		#10 PDB = 24'h12;
		
// 		#10 PDB = 24'h000000;
// 			YDB_in = 24'h133;
		
// 		#10	PDB = 24'b00000101_0_1_110000_0_0_1_00000;	/* m0, x:#56 */
// 			YDB_in = 24'hzzzzzz;

//		#10 PDB = 24'h56;
		

		/* MOVEC Class II */
		/*                     W   aaaaaa   s   ddddd */
// 		#10 PDB = 24'b00000101_0_0_011001_0_0_1_00010;	/* m2, x:#19 */

// 		#10 PDB = 24'h000000;
		
// 		#10 PDB = 24'b00000101_1_0_110011_0_1_1_00100;	/* y:#33, m6 */
		
// 		#10 PDB = 24'h000000;
		
//  	#10 YDB_in = 24'h4141;
//  		PDB = 24'b00000101_0_1_011001_0_0_1_00100;	/* m6, x:(r1)+ */

// 		#10	YDB_in = 24'hzzzzzz;
//  		PDB = 24'h000000;
		


		/* MOVEC Class IV */
		/*                     iiiiiiii     ddddd */
//		#10 PDB = 24'b00000101_00010100_101_00010;	/* #14, m2 */

//		#10 PDB = 24'h000000;
		
//		#10 PDB = 24'b00000101_0_1_011001_0_0_1_00010;	/* m2, x:(r1)+ */


		/* NEG */
		/*                                   d       */
//		#10 PDB = 24'b00000000_00000000_0011_1_110;




		/* REP  Class I  +  NORM */
		/*                        MMMRRR   S        */
//		#10 PDB = 24'b00000110_01_011000_0_0_100000;	/* REP x:(r0)+ */

		/*                           RRR      d      */
//		#10 PDB = 24'b00000001_11011_011_0001_0_101;	/* NORM	R3 <= FFD2 */

//		#10	XDB_in = 24'h2F;
//			PDB = 24'hzzzzzz;

//		#10	XDB_in = 24'h1;
//		    PDB = 24'b001_10111_11111111_00000000; /* I:  r7 = FF */

//		#10 XDB_in = 24'hzzzzzz;		

//		 PDB = 24'b001_10111_11111111_00000000; /* I:  r7 = FF */
			 
//		PDB = 24'h000000;



		/* REP  Class II  +  NORM */
		/*                        aaaaaa   S        */
//		#10 PDB = 24'b00000110_00_010000_0_0_100000;	/* REP x:$10 */

		/*                           RRR      d      */
//		#10 PDB = 24'b00000001_11011_011_0001_0_101;	/* NORM	R3 <= FFD2 */

//		#10	XDB_in = 24'h2f;
//			PDB = 24'hzzzzzz;
		
//		#460 XDB_in = 24'hzzzzzz;
//		 PDB = 24'b001_10111_11111111_00000000; /* I:  r7 = FF */
			 
//		PDB = 24'h000000;



		/* REP  Class III  +  NORM */
		/*                     iiiiiiii      hhhh     */
//		#10 PDB = 24'b00000110_00101111_1010_0000;	/* REP #2F */
//		#10 PDB = 24'b00000110_00000101_1010_0000;	/* REP #5 */
//		#10 PDB = 24'b00000110_00000010_1010_0000;	/* REP #2 */
//		#10 PDB = 24'b00000110_00000011_1010_0000;	/* REP #3 */
//		#10 PDB = 24'b00000110_00000001_1010_0000;	/* REP #1 */

		/*                           RRR      d      */
//		#10 PDB = 24'b00000001_11011_011_0001_0_101;	/* NORM	R3 <= (for #2F rep) FFD2 */

//		#10	PDB = 24'hzzzzzz;

//		#460 PDB = 24'b001_10111_11111111_00000000; /* I:  r7 = FF */

//		#10	PDB = 24'h000000;
		


		/* REP  Class IV  +  NORM */
		/*                                 */
//		#10 PDB = 24'b001_10000_00101111_00000000; /* I: R0 <= #2F */

//		#10	PDB = 24'h000000;

		/*                        dddddd            */
//		#10 PDB = 24'b00000110_11_010000_00100000;	/* REP r0 */

		/*                           RRR      d      */
//		#10 PDB = 24'b00000001_11011_011_0001_0_101;	/* NORM	R3 <= FFD2 */

//		#10	PDB = 24'hzzzzzz;

//		#460 PDB = 24'b001_10111_11111111_00000000; /* I:  r7 = FF */

//		#10	PDB = 24'h000000;



//		#10 PDB = 24'b001_01011_00101111_00000000; /* I: B2 <= #2F */

//		#10	PDB = 24'h000000;

		/*                        dddddd            */
//		#10 PDB = 24'b00000110_11_001011_00100000;	/* REP B2 */

		/*                           RRR      d      */
//		#10 PDB = 24'b00000001_11011_011_0001_0_101;	/* NORM	R3 <= FFD2 */

//		#10	PDB = 24'hzzzzzz;

//		#460 PDB = 24'b001_10111_11111111_00000000; /* I:  r7 = FF */

//		#10	PDB = 24'h000000;




		/* RND */
		/*                                   d      */
//		#10 PDB = 24'b00000000_00000000_0001_0_001;


		/* ROL */
		/*                                   d       */
//		#10 PDB = 24'b00000000_00000000_0011_0_111;


		/* SUB */
		/*                                JJJ d      */
//		#10 PDB = 24'b00000000_00000000_0_110_0_100;


		/* TST */
		/*                                   d      */
//		#10 PDB = 24'b00000000_00000000_0000_0_011;






		#10 PDB = 24'h000000;


		#200 $finish;		/* end simulation */
		
		$shm_close;		/* close the dump file */
	end



/*==============================================================================*/
/*	clock	5 units High, 5 units Low											*/
/*==============================================================================*/

always
	begin
		#5 Clk = 1;
		#5 Clk = 0;
	end
	





endmodule	/* end module top */
